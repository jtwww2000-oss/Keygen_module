`timescale 1ns / 1ps

(* use_dsp48="no" *) // LUT ���ұ���Ҫ���� DSP
module g1_rom(
    g1,
    mid,
    clk
);

    output reg [23:0] g1;
    input      [8:0]  mid;
    input             clk;

    reg [23:0] lut_val;

    // ����߼����ұ�
    always @(*) begin
        case(mid)
            // Mid = 1 (Step 9) -> g^256 mod Q = -1
            9'd1:   lut_val = 24'd8380416; 
            
            // Mid = 2 (Step 8) -> g^128 mod Q
            9'd2:   lut_val = 24'd4808194;   
            
            // Mid = 4 (Step 7) -> g^64 mod Q
            9'd4:   lut_val = 24'd3765607; 
            
            // Mid = 8 (Step 6) -> g^32 mod Q
            9'd8:   lut_val = 24'd5178923;  
            
            // Mid = 16 (Step 5) -> g^16 mod Q
            9'd16:  lut_val = 24'd7778734; 
            
            // Mid = 32 (Step 4) -> g^8 mod Q
            9'd32:  lut_val = 24'd5010068; 
            
            // Mid = 64 (Step 3) -> g^4 mod Q
            9'd64:  lut_val = 24'd3602218; 
            
            // Mid = 128 (Step 2) -> g^2 mod Q
            9'd128: lut_val = 24'd3073009; 
            
            // �쳣������� mid=100 ��������2�ݴ�ֵ��Ĭ�Ϸ��� 1 �򱨴�
            // ��ʵ�� NTT �У������״̬���ܷ���
            default: lut_val = 24'd1;
        endcase
    end

    // ʱ���߼���� (��һ��)
    always @(posedge clk) begin
        g1 <= lut_val;
    end

endmodule