`timescale 1ns / 1ps

module mod_add #(
    parameter WIDTH = 24
)(
    input  wire [WIDTH-1:0] a,
    input  wire [WIDTH-1:0] b,
    input  wire [WIDTH-1:0] q, // Modulus
    output wire [WIDTH-1:0] res
);

    wire [WIDTH:0] sum;
    
    // ���� a + b
    assign sum = a + b;
    
    // ����� >= q�����ȥ q������ֱ�����
    // ����һ��������߼�ѡ����
    assign res = (sum >= q) ? (sum - q) : sum[WIDTH-1:0];

endmodule