`timescale 1ns / 1ps

module Rejsam_a (
    input  wire                 clk,
    input  wire                 rst_n,
    
    // --- ���ƽӿ� ---
    input  wire                 i_start,        // �����ź�
    input  wire [255:0]         i_rho,          // rho (256 bits)
    input  wire [7:0]           i_row,          // ������ row
    input  wire [7:0]           i_column,       // ������ column
    
    // --- ����ӿ� (��ʽ���) ---
    output reg                  o_coeff_valid,  // ϵ����Ч��־
    output reg  [22:0]          o_coeff_data,   // ���ɵ�ϵ�� (< 8380417)
    output reg                  o_done          // ����ź� (������ 256 ��ϵ��)
);

    // --- �������� ---
    localparam Q_VAL = 23'd8380417;
    localparam CNT_TARGET = 9'd256;
    
    // SHAKE128 ����
    localparam RATE_BYTES = 168;            // SHAKE128 Rate = 1344 bits = 168 bytes
    localparam ABSORB_LEN = 256 + 8 + 8;    // rho(256) + col(8) + row(8) = 272 bits

    // --- ״̬�� ---
    localparam S_IDLE        = 3'd0;
    localparam S_START_SHAKE = 3'd1;
    localparam S_REQ_SQUEEZE = 3'd2;
    localparam S_WAIT_DATA   = 3'd3;
    localparam S_PROCESS     = 3'd4;
    localparam S_DONE        = 3'd5;
    // ����״̬���ȴ�����Ӧ��
    localparam S_WAIT_ACK    = 3'd6;

    reg [2:0] state;
    
    // --- �ڲ��ź� ---
    reg [8:0] coeff_cnt;                    // �����ɵ�ϵ������ (0-256)
    reg [10:0] bit_ptr;                     // ��ǰ������ bit ָ�� (0-1344)
    
    // SHAKE128 �ӿ��ź�
    reg  shake_start;
    wire [ABSORB_LEN-1:0] shake_seed;
    wire shake_busy;
    reg  shake_squeeze_req;
    wire shake_squeeze_valid;
    wire [RATE_BYTES*8-1:0] shake_out_data;
    
    // ���� SHAKE ��������ݿ�
    reg [RATE_BYTES*8-1:0] data_buffer;

    // --- 1. �������� Seed ---
    // MATLAB: [rho, column, row] (���� 1 �� LSB)
    // Verilog: {row, column, rho}
    assign shake_seed = {i_row, i_column, i_rho};

    // --- 2. ʵ���� SHAKE128 ---
    // ע�⣺��ȷ����� SHAKE128 ģ���������˴�һ��
    SHAKE128 #(
        .OUTPUT_LEN_BYTES(RATE_BYTES), // ÿ�� Squeeze ��� 168 �ֽ�
        .ABSORB_LEN(ABSORB_LEN)        // ���� 272 bits
    ) u_shake128 (
        .clk             (clk),
        .rst_n           (rst_n),
        .i_start         (shake_start),
        .i_seed          (shake_seed),
        .o_busy          (shake_busy),
        .i_squeeze_req   (shake_squeeze_req),
        .o_squeeze_valid (shake_squeeze_valid),
        .o_squeeze_data  (shake_out_data)
    );

    // --- 3. ���߼� ---
    
    // ��ѡֵ��ȡ (�� buffer ��ȡ 24 bits)
    wire [23:0] raw_chunk;
    wire [22:0] candidate;
    
    // ��̬��Ƭ: ȡ buffer[bit_ptr +: 24]
    // ע��: Verilog ��֧�ֱ�����Ϊ +: ��������ַ��ͨ����Ҫ�� generate �� case��
    // �����������ǿ���ͨ����λ buffer ��ʵ����ʽ����
    // Ϊ�˽�ʡ����������� S_PROCESS ״̬���ƶ� bit_ptr�� combinational logic ��ȡ
    assign raw_chunk = data_buffer[bit_ptr +: 24];
    
    // ��Ӧ MATLAB: bin2dec(flip(...)) ȡ 23 bits
    // ����� raw_chunk[22:0] ��Ϊ�� 23 λ
    assign candidate = raw_chunk[22:0];

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_IDLE;
            o_coeff_valid <= 1'b0;
            o_coeff_data  <= 23'd0;
            o_done <= 1'b0;
            shake_start <= 1'b0;
            shake_squeeze_req <= 1'b0;
            coeff_cnt <= 9'd0;
            bit_ptr <= 11'd0;
            data_buffer <= 0;
        end else begin
            // Ĭ�����帴λ
            shake_start <= 1'b0;
            shake_squeeze_req <= 1'b0;
            o_coeff_valid <= 1'b0; // valid �ź�ֻά��һ��

            case (state)
                S_IDLE: begin
                    o_done <= 1'b0;
                    coeff_cnt <= 9'd0;
                    if (i_start) begin
                        state <= S_START_SHAKE;
                    end
                end

                S_START_SHAKE: begin
                    shake_start <= 1'b1; // ���� SHAKE ����
                    state <= S_REQ_SQUEEZE; // ֱ��ȥ������� (One-Shot ģʽ���Զ����� absorb)
                end

                S_REQ_SQUEEZE: begin
                    // �ȴ� SHAKE æ�����գ�����æ����һ�� squeeze
                    // ע�⣺����֮ǰ����ƣ�busy Ϊ 1 ʱ���ܲ�������ȴ� busy ����ٱ�ͣ�
                    // ֮ǰ�� SHAKE Controller ����ǣ�Start -> Busy=1 -> Valid -> SqueezeReq -> Valid...
                    // �������ǵȴ� shake_busy ���(������Ѿ��������) ����ֱ�ӿ� squeeze_valid
                    // Ϊ���Ƚ������Ƿ�������
                    // ���� SHAKE ģ���� absorb ��ɺ���Զ����� SQUEEZE ״̬���ȴ� req
                    shake_squeeze_req <= 1'b1;
                    state <= S_WAIT_ACK;
                end
                
                
                S_WAIT_ACK: begin
                    shake_squeeze_req <= 1'b0; // ������������
                    
                    // ������ͣһ�ģ��� SHAKE ģ��ʱ��ȥ��Ӧ req ���� valid ����
                    // ����������һ��״̬ʱ��valid �ͻ����ȵ��� 0 ��
                    if (shake_squeeze_valid == 1'b0) begin
                         state <= S_WAIT_DATA;
                    end
                    // ��� SHAKE ��Ӧ����valid ��û��ͣ�����������������
                    // (ͨ��һ�ľ͹���ֱ�� else state <= S_WAIT_DATA Ҳ���ԣ������жϸ��Ƚ�)
                end
                
                
                S_WAIT_DATA: begin
                    if (shake_squeeze_valid) begin
                        data_buffer <= shake_out_data;
                        bit_ptr <= 11'd0; // ����ָ�뵽 buffer ͷ�� (LSB)
                        state <= S_PROCESS;
                    end
                end

                S_PROCESS: begin
                    // ����Ƿ� buffer ʣ�಻�� 24 bits
                    // 1344 - 24 = 1320. ��� ptr > 1320��˵��ʣ�µĲ�����
                    if (bit_ptr > (RATE_BYTES*8 - 24)) begin
                        // Buffer �����ˣ���Ҫ��������
                        state <= S_REQ_SQUEEZE;
                    end else begin
                        // ��鵱ǰ��ѡֵ
                        if (candidate < Q_VAL) begin
                            o_coeff_valid <= 1'b1;
                            o_coeff_data <= candidate;
                            coeff_cnt <= coeff_cnt + 1;
                            
                            // ����Ƿ����
                            if (coeff_cnt == (CNT_TARGET - 1)) begin
                                state <= S_DONE;
                            end
                        end
                        
                        // �ƶ�ָ�� (������һ�� 24 bits)
                        // ��Ӧ MATLAB: ѭ�� i �� 1��ÿ������ 24 bits
                        bit_ptr <= bit_ptr + 24; 
                    end
                end

                S_DONE: begin
                    o_done <= 1'b1;
                    // �ȴ��ⲿ��λ���µ� start
                    if (i_start) begin
                        state <= S_START_SHAKE;
                        o_done <= 1'b0;
                        coeff_cnt <= 9'd0;
                    end
                end
            endcase
        end
    end

endmodule