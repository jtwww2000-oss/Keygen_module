`timescale 1ns / 1ps

module Barrett_reduce #(
    parameter WIDTH = 24
)(
    input  wire               clk,
    input  wire [2*WIDTH-1:0] prod, // ����˻� (48 bits)
    input  wire [WIDTH-1:0]   q,    // Modulus Q
    input  wire [WIDTH+1:0]   mu,   // Constant mu (2^48 / Q)
    output reg  [WIDTH-1:0]   res
);

    // --------------------------------------------------------
    // Stage 1: �����̵ĵ�һ�� big_prod = prod * mu
    // --------------------------------------------------------
    (* use_dsp = "yes" *) reg [3*WIDTH+1:0] r1_big_prod;
    reg [2*WIDTH-1:0] r1_prod; // ����ԭʼ����
    reg [WIDTH-1:0]   r1_q;

    always @(posedge clk) begin
        r1_big_prod <= prod * mu;
        r1_prod     <= prod;
        r1_q        <= q;
    end

    // --------------------------------------------------------
    // Stage 2: ������� sub_term = floor(...) * q
    // --------------------------------------------------------
    (* use_dsp = "yes" *) reg [WIDTH+2:0] r2_q_times_qhat;
    reg [WIDTH+2:0]   r2_prod_low; // ֻ��Ҫ������λ���ڼ���
    reg [WIDTH-1:0]   r2_q;

    wire [WIDTH+2:0] q_hat;
    
    // ���� �����㣺�������� 48 λ (ƥ�� mu = 2^48 / Q) ����
    assign q_hat = r1_big_prod >> 48; 

    always @(posedge clk) begin
        r2_q_times_qhat <= q_hat * r1_q;
        // ����ֻ��Ҫ prod �ĵ�λ���������ļ����Ƚ�
        // ȡ 27 λ�㹻���ɲ��� (WIDTH + 3)
        r2_prod_low     <= r1_prod[WIDTH+2:0]; 
        r2_q            <= r1_q;
    end

    // --------------------------------------------------------
    // Stage 3: ���ռ���������
    // --------------------------------------------------------
    wire [WIDTH+2:0] r_raw;
    wire [WIDTH+2:0] r_corr;
    wire [WIDTH-1:0] r_final;

    assign r_raw = r2_prod_low - r2_q_times_qhat;
    
    // �����߼�
    assign r_corr  = (r_raw >= r2_q) ? (r_raw - r2_q) : r_raw;
    assign r_final = (r_corr >= r2_q) ? (r_corr - r2_q) : r_corr[WIDTH-1:0];

    always @(posedge clk) begin
        res <= r_final;
    end

endmodule