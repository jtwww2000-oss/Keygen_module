//`timescale 1ns / 1ps

//module pad #(
//    parameter X = 1088,          // Rate (SHAKE256)
//    parameter MAX_LEN = 1088     // ��������С
//)(
//    input  wire [MAX_LEN-1:0]        N,     // ������Ϣ���� N (��λ����)
//    input  wire [$clog2(MAX_LEN)-1:0] m,     // ������Ϣ���� (bits)
//    output reg  [MAX_LEN-1:0]        P      // ��� P
//);

//    // ���� SHAKE256 ��ָ��� (4 bits)
//    // ע�⣺���ﶨ��Ϊ 4'b1111��
//    // ������ MATLAB �Ǹ�λ�ں���߼����� 4 λ�ᱻ�ŵ� N �ĸ�λ����
//    localparam [3:0] DOMAIN_SEP = 4'b1111;

//    integer i;

//    always @(*) begin
//        // 1. ��ʼ�� P Ϊȫ 0
//        // ��һ���ǳ���Ҫ�����Զ�������м�� 0 (j��0)
//        P = {MAX_LEN{1'b0}};

//        // 2. �������� N
//        // N �������λ [0 �� m-1]
//        // Ϊ���ۺ����Ѻã�����ʹ�ü򵥵������߼���ֱ�Ӹ�ֵ
//        // (ע�⣺������������ N �� m λ���ϱ������ 0��������ǣ���Ҫ�ض�)
//        // �ڷ����߼��У����ͬ��: P[m-1:0] = N[m-1:0];
//        // �� Verilog ��֧�ֱ�����Χ��Ƭ����������ֱ��ȫ��ֵ�������������ǻ���� N ��λ����
//        P = N; 

//        // 3. ���� SHAKE256 ��ָ��� '1111'
//        // λ�ã����������� N �ĸ�λ����
//        // ������Χ��[m+3 : m]
//        // ����ȫ���� "1111 �� N �ĸ�λ" ��һ����
//        for (i = 0; i < 4; i = i + 1) begin
//            P[m + i] = DOMAIN_SEP[i];
//        end
        
//        // 4. ���� Padding Start '1'
//        // λ�ã�����ָ�������һλ
//        // ������m + 4
//        P[m + 4] = 1'b1;

//        // 5. ���� Padding End '1'
//        // λ�ã�Rate �����λ (X-1)
//        // ��Ӧ MATLAB P �����һ��Ԫ��
//        P[X - 1] = 1'b1;
        
//        // ���䣺�����ص� (Overlap)
//        // ��� m + 4 �պõ��� X - 1 (��������÷ǳ���)��
//        // ����ĸ�ֵ���Ⱥ��ͬһ�� bit ���в�����
//        // ��Ϊ������ 1�������߼����Ǽ��ݵ� (1 | 1 = 1)��
//        // ��Ϊ���Ͻ���Verilog ��������ֵ '=' ��һ���Ḳ��ǰһ����
//        // ��Ϊ P[X-1] = 1 �����ִ�еģ���������������λ���� 1������ Sponge �淶��
//    end

//endmodule


`timescale 1ns / 1ps
module pad #(
    parameter X = 1088,          // Rate
    parameter MAX_LEN = 1088     // Buffer Size
)(
    input  wire [MAX_LEN-1:0]        N,
    input  wire [$clog2(MAX_LEN)-1:0] m,
    output reg  [MAX_LEN-1:0]        P
);

    localparam [3:0] DOMAIN_SEP = 4'b1111;

    always @(*) begin
        // 1. �ȸ������� (���� N ��λ�Ѳ�0)
        P = N; 
        
        // 2. ���� SHAKE256 ��ָ��� '1111'
        // ʹ�� Verilog-2001 "Indexed Part Select" �﷨: [base +: width]
        // �� m ��ʼ������ȡ 4 λ
        P[m +: 4] = DOMAIN_SEP;
        
        // 3. ���� Padding Start '1'
        // ע�⣺m+4 �ǽ�������ָ�������һλ
        P[m + 4] = 1'b1;
        
        // 4. ���� Padding End '1' at Rate block boundary
        P[X - 1] = 1'b1;
    end

endmodule